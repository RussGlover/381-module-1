package fft_len is
constant LOG2_FFT_LEN : integer := 10;
end fft_len;